
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mem is
port(
    addr: std_ulogic_vector(7 downto 0);
    dout: out std_ulogic_vector(31 downto 0) := (others => '0'));
end entity;


architecture impl of mem is
    type mem_t is array(natural range 0 to 255) of
        std_ulogic_vector(31 downto 0);
    constant data: mem_t := (

        std_ulogic_vector(to_unsigned(4852, 32)),
        std_ulogic_vector(to_unsigned(4938, 32)),
        std_ulogic_vector(to_unsigned(5625, 32)),
        std_ulogic_vector(to_unsigned(6260, 32)),
        std_ulogic_vector(to_unsigned(1904, 32)),
        std_ulogic_vector(to_unsigned(76  , 32)),
        std_ulogic_vector(to_unsigned(8245, 32)),
        std_ulogic_vector(to_unsigned(1231, 32)),
        std_ulogic_vector(to_unsigned(7294, 32)),
        std_ulogic_vector(to_unsigned(6598, 32)),
        std_ulogic_vector(to_unsigned(7457, 32)),
        std_ulogic_vector(to_unsigned(5769, 32)),
        std_ulogic_vector(to_unsigned(4171, 32)),
        std_ulogic_vector(to_unsigned(7690, 32)),
        std_ulogic_vector(to_unsigned(5970, 32)),
        std_ulogic_vector(to_unsigned(3615, 32)),
        std_ulogic_vector(to_unsigned(6246, 32)),
        std_ulogic_vector(to_unsigned(6695, 32)),
        std_ulogic_vector(to_unsigned(4825, 32)),
        std_ulogic_vector(to_unsigned(5217, 32)),
        std_ulogic_vector(to_unsigned(9495, 32)),
        std_ulogic_vector(to_unsigned(8642, 32)),
        std_ulogic_vector(to_unsigned(7611, 32)),
        std_ulogic_vector(to_unsigned(8862, 32)),
        std_ulogic_vector(to_unsigned(5248, 32)),
        std_ulogic_vector(to_unsigned(1397, 32)),
        std_ulogic_vector(to_unsigned(87  , 32)),
        std_ulogic_vector(to_unsigned(4431, 32)),
        std_ulogic_vector(to_unsigned(1333, 32)),
        std_ulogic_vector(to_unsigned(8134, 32)),
        std_ulogic_vector(to_unsigned(8882, 32)),
        std_ulogic_vector(to_unsigned(1870, 32)),
        std_ulogic_vector(to_unsigned(6265, 32)),
        std_ulogic_vector(to_unsigned(9539, 32)),
        std_ulogic_vector(to_unsigned(9444, 32)),
        std_ulogic_vector(to_unsigned(3040, 32)),
        std_ulogic_vector(to_unsigned(3656, 32)),
        std_ulogic_vector(to_unsigned(7956, 32)),
        std_ulogic_vector(to_unsigned(1380, 32)),
        std_ulogic_vector(to_unsigned(6048, 32)),
        std_ulogic_vector(to_unsigned(6525, 32)),
        std_ulogic_vector(to_unsigned(1100, 32)),
        std_ulogic_vector(to_unsigned(1198, 32)),
        std_ulogic_vector(to_unsigned(1525, 32)),
        std_ulogic_vector(to_unsigned(7604, 32)),
        std_ulogic_vector(to_unsigned(2415, 32)),
        std_ulogic_vector(to_unsigned(946 , 32)),
        std_ulogic_vector(to_unsigned(8541, 32)),
        std_ulogic_vector(to_unsigned(9730, 32)),
        std_ulogic_vector(to_unsigned(7322, 32)),
        std_ulogic_vector(to_unsigned(1581, 32)),
        std_ulogic_vector(to_unsigned(8978, 32)),
        std_ulogic_vector(to_unsigned(5484, 32)),
        std_ulogic_vector(to_unsigned(6669, 32)),
        std_ulogic_vector(to_unsigned(5568, 32)),
        std_ulogic_vector(to_unsigned(3549, 32)),
        std_ulogic_vector(to_unsigned(5960, 32)),
        std_ulogic_vector(to_unsigned(6834, 32)),
        std_ulogic_vector(to_unsigned(7503, 32)),
        std_ulogic_vector(to_unsigned(2874, 32)),
        std_ulogic_vector(to_unsigned(8347, 32)),
        std_ulogic_vector(to_unsigned(8437, 32)),
        std_ulogic_vector(to_unsigned(6641, 32)),
        std_ulogic_vector(to_unsigned(5218, 32)),
        std_ulogic_vector(to_unsigned(1115, 32)),
        std_ulogic_vector(to_unsigned(5262, 32)),
        std_ulogic_vector(to_unsigned(8196, 32)),
        std_ulogic_vector(to_unsigned(9183, 32)),
        std_ulogic_vector(to_unsigned(2459, 32)),
        std_ulogic_vector(to_unsigned(592 , 32)),
        std_ulogic_vector(to_unsigned(972 , 32)),
        std_ulogic_vector(to_unsigned(1882, 32)),
        std_ulogic_vector(to_unsigned(7456, 32)),
        std_ulogic_vector(to_unsigned(366 , 32)),
        std_ulogic_vector(to_unsigned(1883, 32)),
        std_ulogic_vector(to_unsigned(2682, 32)),
        std_ulogic_vector(to_unsigned(2697, 32)),
        std_ulogic_vector(to_unsigned(379 , 32)),
        std_ulogic_vector(to_unsigned(8497, 32)),
        std_ulogic_vector(to_unsigned(6127, 32)),
        std_ulogic_vector(to_unsigned(4397, 32)),
        std_ulogic_vector(to_unsigned(8773, 32)),
        std_ulogic_vector(to_unsigned(8645, 32)),
        std_ulogic_vector(to_unsigned(17  , 32)),
        std_ulogic_vector(to_unsigned(383 , 32)),
        std_ulogic_vector(to_unsigned(6968, 32)),
        std_ulogic_vector(to_unsigned(7458, 32)),
        std_ulogic_vector(to_unsigned(4893, 32)),
        std_ulogic_vector(to_unsigned(4907, 32)),
        std_ulogic_vector(to_unsigned(4798, 32)),
        std_ulogic_vector(to_unsigned(641 , 32)),
        std_ulogic_vector(to_unsigned(4042, 32)),
        std_ulogic_vector(to_unsigned(5746, 32)),
        std_ulogic_vector(to_unsigned(1500, 32)),
        std_ulogic_vector(to_unsigned(9456, 32)),
        std_ulogic_vector(to_unsigned(903 , 32)),
        std_ulogic_vector(to_unsigned(1922, 32)),
        std_ulogic_vector(to_unsigned(5293, 32)),
        std_ulogic_vector(to_unsigned(617 , 32)),
        std_ulogic_vector(to_unsigned(4674, 32)),
        std_ulogic_vector(to_unsigned(2482, 32)),
        std_ulogic_vector(to_unsigned(9752, 32)),
        std_ulogic_vector(to_unsigned(1131, 32)),
        std_ulogic_vector(to_unsigned(5867, 32)),
        std_ulogic_vector(to_unsigned(4945, 32)),
        std_ulogic_vector(to_unsigned(2446, 32)),
        std_ulogic_vector(to_unsigned(387 , 32)),
        std_ulogic_vector(to_unsigned(5831, 32)),
        std_ulogic_vector(to_unsigned(7522, 32)),
        std_ulogic_vector(to_unsigned(5828, 32)),
        std_ulogic_vector(to_unsigned(3440, 32)),
        std_ulogic_vector(to_unsigned(3255, 32)),
        std_ulogic_vector(to_unsigned(8232, 32)),
        std_ulogic_vector(to_unsigned(5035, 32)),
        std_ulogic_vector(to_unsigned(4970, 32)),
        std_ulogic_vector(to_unsigned(9264, 32)),
        std_ulogic_vector(to_unsigned(2425, 32)),
        std_ulogic_vector(to_unsigned(1884, 32)),
        std_ulogic_vector(to_unsigned(6718, 32)),
        std_ulogic_vector(to_unsigned(6884, 32)),
        std_ulogic_vector(to_unsigned(1026, 32)),
        std_ulogic_vector(to_unsigned(9204, 32)),
        std_ulogic_vector(to_unsigned(4177, 32)),
        std_ulogic_vector(to_unsigned(2381, 32)),
        std_ulogic_vector(to_unsigned(6500, 32)),
        std_ulogic_vector(to_unsigned(6825, 32)),
        std_ulogic_vector(to_unsigned(6305, 32)),
        std_ulogic_vector(to_unsigned(4577, 32)),
        std_ulogic_vector(to_unsigned(8001, 32)),
        std_ulogic_vector(to_unsigned(3410, 32)),
        std_ulogic_vector(to_unsigned(5088, 32)),
        std_ulogic_vector(to_unsigned(6609, 32)),
        std_ulogic_vector(to_unsigned(8081, 32)),
        std_ulogic_vector(to_unsigned(2672, 32)),
        std_ulogic_vector(to_unsigned(2956, 32)),
        std_ulogic_vector(to_unsigned(4189, 32)),
        std_ulogic_vector(to_unsigned(4384, 32)),
        std_ulogic_vector(to_unsigned(5875, 32)),
        std_ulogic_vector(to_unsigned(2919, 32)),
        std_ulogic_vector(to_unsigned(7376, 32)),
        std_ulogic_vector(to_unsigned(6521, 32)),
        std_ulogic_vector(to_unsigned(8311, 32)),
        std_ulogic_vector(to_unsigned(9912, 32)),
        std_ulogic_vector(to_unsigned(6528, 32)),
        std_ulogic_vector(to_unsigned(2320, 32)),
        std_ulogic_vector(to_unsigned(6098, 32)),
        std_ulogic_vector(to_unsigned(9521, 32)),
        std_ulogic_vector(to_unsigned(8374, 32)),
        std_ulogic_vector(to_unsigned(3215, 32)),
        std_ulogic_vector(to_unsigned(1707, 32)),
        std_ulogic_vector(to_unsigned(7174, 32)),
        std_ulogic_vector(to_unsigned(6064, 32)),
        std_ulogic_vector(to_unsigned(423 , 32)),
        std_ulogic_vector(to_unsigned(7493, 32)),
        std_ulogic_vector(to_unsigned(4294, 32)),
        std_ulogic_vector(to_unsigned(6705, 32)),
        std_ulogic_vector(to_unsigned(9788, 32)),
        std_ulogic_vector(to_unsigned(8531, 32)),
        std_ulogic_vector(to_unsigned(5999, 32)),
        std_ulogic_vector(to_unsigned(567 , 32)),
        std_ulogic_vector(to_unsigned(1328, 32)),
        std_ulogic_vector(to_unsigned(2430, 32)),
        std_ulogic_vector(to_unsigned(7424, 32)),
        std_ulogic_vector(to_unsigned(2276, 32)),
        std_ulogic_vector(to_unsigned(159 , 32)),
        std_ulogic_vector(to_unsigned(9292, 32)),
        std_ulogic_vector(to_unsigned(4812, 32)),
        std_ulogic_vector(to_unsigned(5801, 32)),
        std_ulogic_vector(to_unsigned(9799, 32)),
        std_ulogic_vector(to_unsigned(3211, 32)),
        std_ulogic_vector(to_unsigned(261 , 32)),
        std_ulogic_vector(to_unsigned(7878, 32)),
        std_ulogic_vector(to_unsigned(7753, 32)),
        std_ulogic_vector(to_unsigned(698 , 32)),
        std_ulogic_vector(to_unsigned(3056, 32)),
        std_ulogic_vector(to_unsigned(2217, 32)),
        std_ulogic_vector(to_unsigned(9404, 32)),
        std_ulogic_vector(to_unsigned(466 , 32)),
        std_ulogic_vector(to_unsigned(7209, 32)),
        std_ulogic_vector(to_unsigned(3373, 32)),
        std_ulogic_vector(to_unsigned(1476, 32)),
        std_ulogic_vector(to_unsigned(9669, 32)),
        std_ulogic_vector(to_unsigned(177 , 32)),
        std_ulogic_vector(to_unsigned(7026, 32)),
        std_ulogic_vector(to_unsigned(4689, 32)),
        std_ulogic_vector(to_unsigned(1534, 32)),
        std_ulogic_vector(to_unsigned(7227, 32)),
        std_ulogic_vector(to_unsigned(3324, 32)),
        std_ulogic_vector(to_unsigned(1851, 32)),
        std_ulogic_vector(to_unsigned(3425, 32)),
        std_ulogic_vector(to_unsigned(190 , 32)),
        std_ulogic_vector(to_unsigned(3196, 32)),
        std_ulogic_vector(to_unsigned(919 , 32)),
        std_ulogic_vector(to_unsigned(2332, 32)),
        std_ulogic_vector(to_unsigned(6397, 32)),
        std_ulogic_vector(to_unsigned(7965, 32)),
        std_ulogic_vector(to_unsigned(8658, 32)),
        std_ulogic_vector(to_unsigned(2988, 32)),
        std_ulogic_vector(to_unsigned(2984, 32)),
        std_ulogic_vector(to_unsigned(6946, 32)),
        std_ulogic_vector(to_unsigned(9083, 32)),
        std_ulogic_vector(to_unsigned(1873, 32)),
        std_ulogic_vector(to_unsigned(9330, 32)),
        std_ulogic_vector(to_unsigned(6980, 32)),
        std_ulogic_vector(to_unsigned(5201, 32)),
        std_ulogic_vector(to_unsigned(4305, 32)),
        std_ulogic_vector(to_unsigned(2503, 32)),
        std_ulogic_vector(to_unsigned(864 , 32)),
        std_ulogic_vector(to_unsigned(945 , 32)),
        std_ulogic_vector(to_unsigned(7454, 32)),
        std_ulogic_vector(to_unsigned(2060, 32)),
        std_ulogic_vector(to_unsigned(9349, 32)),
        std_ulogic_vector(to_unsigned(8750, 32)),
        std_ulogic_vector(to_unsigned(7968, 32)),
        std_ulogic_vector(to_unsigned(6574, 32)),
        std_ulogic_vector(to_unsigned(4705, 32)),
        std_ulogic_vector(to_unsigned(3627, 32)),
        std_ulogic_vector(to_unsigned(6063, 32)),
        std_ulogic_vector(to_unsigned(324 , 32)),
        std_ulogic_vector(to_unsigned(4816, 32)),
        std_ulogic_vector(to_unsigned(5338, 32)),
        std_ulogic_vector(to_unsigned(6295, 32)),
        std_ulogic_vector(to_unsigned(679 , 32)),
        std_ulogic_vector(to_unsigned(65  , 32)),
        std_ulogic_vector(to_unsigned(4589, 32)),
        std_ulogic_vector(to_unsigned(3308, 32)),
        std_ulogic_vector(to_unsigned(3989, 32)),
        std_ulogic_vector(to_unsigned(7024, 32)),
        std_ulogic_vector(to_unsigned(7167, 32)),
        std_ulogic_vector(to_unsigned(533 , 32)),
        std_ulogic_vector(to_unsigned(8096, 32)),
        std_ulogic_vector(to_unsigned(4062, 32)),
        std_ulogic_vector(to_unsigned(3904, 32)),
        std_ulogic_vector(to_unsigned(983 , 32)),
        std_ulogic_vector(to_unsigned(7003, 32)),
        std_ulogic_vector(to_unsigned(8570, 32)),
        std_ulogic_vector(to_unsigned(6396, 32)),
        std_ulogic_vector(to_unsigned(7518, 32)),
        std_ulogic_vector(to_unsigned(9484, 32)),
        std_ulogic_vector(to_unsigned(1463, 32)),
        std_ulogic_vector(to_unsigned(7538, 32)),
        std_ulogic_vector(to_unsigned(4929, 32)),
        std_ulogic_vector(to_unsigned(1967, 32)),
        std_ulogic_vector(to_unsigned(6327, 32)),
        std_ulogic_vector(to_unsigned(4360, 32)),
        std_ulogic_vector(to_unsigned(3110, 32)),
        std_ulogic_vector(to_unsigned(8168, 32)),
        std_ulogic_vector(to_unsigned( 907, 32)),
        std_ulogic_vector(to_unsigned( 964, 32)),
        std_ulogic_vector(to_unsigned(9861, 32)),
        std_ulogic_vector(to_unsigned(3075, 32)),
        std_ulogic_vector(to_unsigned(9284, 32)),
        std_ulogic_vector(to_unsigned(2361, 32)),
        std_ulogic_vector(to_unsigned(1389, 32)),
        std_ulogic_vector(to_unsigned(2461, 32)),
        std_ulogic_vector(to_unsigned(9255, 32))

    );
begin

dout <= data(to_integer(unsigned(addr)));

end architecture;
